// dummy dijkstra на всякий пожарный 